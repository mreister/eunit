module counter #( parameter BUS_WIDTH=32)
(
  input logic clock,
  input logic reset,
  output logic [WIDTH-1:0] count
);


end module; 