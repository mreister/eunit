module counter
(
  input logic clock,
  input logic reset,
  output logic [WIDTH-1:0] count
);


end module;